`default_nettype none
// uses 2 BRAMs
module key_schedule (
	input  wire clk,
	input  wire [ 1:0] column,
	input  wire [ 3:0] round,
	output wire [31:0] key // just a column of the state matrix
);

	/*
		iCE40 BRAM fetches two bytes at a time, so to get the
		whole column at once, we need two blocks, one for the
		high bytes and one for the low bytes. Here's the
		human-readable key schedule:

		row       0            1            2            3
		 0   00 01 02 03  04 05 06 07  08 09 0a 0b  0c 0d 0e 0f
		 1   d6 aa 74 fd  d2 af 72 fa  da a6 78 f1  d6 ab 76 fe
		 2   b6 92 cf 0b  64 3d bd f1  be 9b c5 00  68 30 b3 fe
		 3   b6 ff 74 4e  d2 c2 c9 bf  6c 59 0c bf  04 69 bf 41
		 4   47 f7 f7 bc  95 35 3e 03  f9 6c 32 bc  fd 05 8d fd
		 5   3c aa a3 e8  a9 9f 9d eb  50 f3 af 57  ad f6 22 aa
		 6   5e 39 0f 7d  f7 a6 92 96  a7 55 3d c1  0a a3 1f 6b
		 7   14 f9 70 1a  e3 5f e2 8c  44 0a df 4d  4e a9 c0 26
		 8   47 43 87 35  a4 1c 65 b9  e0 16 ba f4  ae bf 7a d2
		 9   54 99 32 d1  f0 85 57 68  10 93 ed 9c  be 2c 97 4e
		 a   13 11 1d 7f  e3 94 4a 17  f3 07 a7 8b  4d 2b 30 c5

		In this view, "round" chooses the row, and "column"
		chooses the set of four bytes within that row.
	*/

	/* ---------------------------------------------- */
	/* === T-tables auto-generated by gen_bram.py === */
	/* ---------------------------------------------- */

	SB_RAM40_4K #(
		.INIT_0(256'h6904596cc2d2ffb630689bbe3d6492b6abd6a6daafd2aad60d0c090805040100),
		.INIT_1(256'ha94e0a445fe3f914a30a55a7a6f7395ef6adf3509fa9aa3c05fd6cf93595f747),
		.INIT_2(256'h00000000000000002b4d07f394e311132cbe931085f09954bfae16e01ca44347)
	) keys_lo (
		.RADDR({5'b0, round, column}),
		.RDATA({key[15:0]}),
		.RCLK (clk),
		.RE   (1'b1),
		.RCLKE(1'b1),
		.WADDR(11'b0),
		.WCLK (1'b0),
		.WCLKE(1'b0),
		.WE   (1'b0),
		.WDATA(16'b0),
		.MASK (16'b0)
	);

	SB_RAM40_4K #(
		.INIT_0(256'h41bfbf0cbfc94e74feb300c5f1bd0bcffe76f178fa72fd740f0e0b0a07060302),
		.INIT_1(256'h26c04ddf8ce21a706b1fc13d96927d0faa2257afeb9de8a3fd8dbc32033ebcf7),
		.INIT_2(256'h0000000000000000c5308ba7174a7f1d4e979ced6857d132d27af4bab9653587)
	) keys_hi (
		.RADDR({5'b0, round, column}),
		.RDATA({key[31:16]}),
		.RCLK (clk),
		.RE   (1'b1),
		.RCLKE(1'b1),
		.WADDR(11'b0),
		.WCLK (1'b0),
		.WCLKE(1'b0),
		.WE   (1'b0),
		.WDATA(16'b0),
		.MASK (16'b0)
	);

endmodule
